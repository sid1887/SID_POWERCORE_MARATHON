module comparator_2bit(
    input wire [1:0] A,B,
    output wire A_gt_B, A_lt_B, A_eq_B
);

assign A_gt_B = (A > B);
assign A_lt_B = (A < B);
assign A_eq_B = (A == B);

endmodule
